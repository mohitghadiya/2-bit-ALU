<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0.763577,-54.582,59.7635,-116.252</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>32,-19.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>32,-23.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AI_XOR2</type>
<position>58,-21</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>71.5,-243.5</position>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_XOR2</type>
<position>72.5,-256</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>51.5,-32.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>74.5,-266</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>43.5,-33.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AI_XOR2</type>
<position>52.5,-45</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>54.5,-55</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>46.5,-56</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AI_XOR2</type>
<position>78,-41</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>89,-49</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AE_SMALL_INVERTER</type>
<position>81.5,-48</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AI_XOR2</type>
<position>98,-252</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR2</type>
<position>96.5,-55</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>109,-260</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>43,-32.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>96.5,-22.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>46.5,-55.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>32.5,-42.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>81,-47.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>31.5,-46</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>116.5,-265.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>102,-41</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>105.5,-54.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>58,-20.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>58,-9.5</position>
<gparam>LABEL_TEXT 2 bit Substraction</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>52,-254.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>29,-20</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>29,-23</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>29.5,-43</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>29,-46.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>100,-22</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>105.5,-40.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>109.5,-54.5</position>
<gparam>LABEL_TEXT Bout</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>23.5,-93</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>23.5,-96</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AI_XOR2</type>
<position>62.5,-94</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>47,-117.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>52,-257.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AI_XOR2</type>
<position>72.5,-103</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>71,-127</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>122,-252</position>
<input>
<ID>N_in0</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AI_XOR2</type>
<position>101,-104</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>98,-116.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>125.5,-265.5</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AE_OR2</type>
<position>105.5,-125.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>GA_LED</type>
<position>116.5,-94.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>46,-101</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>46,-104</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>122.5,-104</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>122,-125.5</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>72,-85.5</position>
<gparam>LABEL_TEXT 2 bit Addition</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>20,-92.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>20.5,-96</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>43,-100.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>43,-103.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>119,-93.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>125.5,-103.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>126,-125</position>
<gparam>LABEL_TEXT Bout</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>160,-24</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>52.5,-44.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>64</ID>
<type>AI_XOR2</type>
<position>177.5,-26.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>179.5,-36.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_SMALL_INVERTER</type>
<position>171.5,-37.5</position>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>67</ID>
<type>AI_XOR2</type>
<position>180.5,-49</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>182.5,-59</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_SMALL_INVERTER</type>
<position>174.5,-60</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AI_XOR2</type>
<position>206,-45</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_AND2</type>
<position>217,-53</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_SMALL_INVERTER</type>
<position>209.5,-52</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR2</type>
<position>224.5,-58.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>224.5,-26.5</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>160,-47.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>230,-45</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>233.5,-58.5</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>157,-24</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>49,-253.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>157.5,-47</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>49.5,-257.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>228,-26</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>233.5,-44.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>237.5,-58.5</position>
<gparam>LABEL_TEXT Bout</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>125.5,-251.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>129.5,-265.5</position>
<gparam>LABEL_TEXT Bout</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>EE_VDD</type>
<position>156,-28.5</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>78,-40.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>91</ID>
<type>FF_GND</type>
<position>159,-51.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>183.5,-15</position>
<gparam>LABEL_TEXT Decrement</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>164,-87</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>164,-90.5</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>AI_XOR2</type>
<position>181.5,-89.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND2</type>
<position>183.5,-99.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AI_XOR2</type>
<position>184.5,-112</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND2</type>
<position>186.5,-122</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AI_XOR2</type>
<position>210,-108</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND2</type>
<position>221,-116</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_OR2</type>
<position>228.5,-121.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>GA_LED</type>
<position>228.5,-89.5</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>164,-110.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>164,-113.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>105</ID>
<type>GA_LED</type>
<position>234,-108</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>GA_LED</type>
<position>237.5,-121.5</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>190.5,-79.5</position>
<gparam>LABEL_TEXT Increment</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>161,-87</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>161,-90</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>161.5,-110</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>161.5,-113.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>232,-89</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>237.5,-107.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>241.5,-121.5</position>
<gparam>LABEL_TEXT Bout</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>51.5,-32</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>54,-54.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_LABEL</type>
<position>88.5,-48.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>96.5,-54.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>62.5,-93.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>72.5,-102.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>46.5,-117</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>98,-116</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>101,-103.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>71,-126.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>105.5,-125</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-20,55,-20</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>34 9</intersection>
<intersection>40 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-33.5,40,-20</points>
<intersection>-33.5 4</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>40,-33.5,41.5,-33.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>40 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>34,-20,34,-19.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-22,55,-22</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>34 7</intersection>
<intersection>42.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-31.5,42.5,-22</points>
<intersection>-31.5 4</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-31.5,48.5,-31.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>42.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>34,-23.5,34,-22</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-33.5,48.5,-33.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-46,49.5,-46</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>45.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45.5,-54,45.5,-46</points>
<intersection>-54 4</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45.5,-54,51.5,-54</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>45.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-56,51.5,-56</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-21,95.5,-21</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>95.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>95.5,-22.5,95.5,-21</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-56,41.5,-42.5</points>
<intersection>-56 4</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-42.5,49.5,-42.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>41.5 0</intersection>
<intersection>49.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-56,44.5,-56</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>49.5,-44,49.5,-42.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-45,65.5,-40</points>
<intersection>-45 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-40,75,-40</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection>
<intersection>69 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-45,65.5,-45</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>65.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69,-48,69,-40</points>
<intersection>-48 4</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>69,-48,79.5,-48</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>69 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-56,75,-55</points>
<intersection>-56 1</intersection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-56,93.5,-56</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-55,75,-55</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-48,86,-48</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-257.5,69.5,-257.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>65.5 3</intersection>
<intersection>69.5 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65.5,-265,65.5,-257.5</points>
<intersection>-265 4</intersection>
<intersection>-257.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>65.5,-265,71.5,-265</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>69.5,-257.5,69.5,-257</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-257.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-41,101,-41</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>25</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-50,25.5,-36.5</points>
<intersection>-50 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-50,86,-50</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection>
<intersection>73 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-36.5,54.5,-36.5</points>
<intersection>25.5 0</intersection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-36.5,54.5,-32.5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>73,-50,73,-42</points>
<intersection>-50 1</intersection>
<intersection>-42 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>73,-42,75,-42</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>73 4</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-54,93,-49</points>
<intersection>-54 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-54,93.5,-54</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,-49,93,-49</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-55,104.5,-55</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>104.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>104.5,-55,104.5,-54.5</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-93,59.5,-93</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>33 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>33,-118.5,33,-93</points>
<intersection>-118.5 6</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>33,-118.5,44,-118.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>33 5</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-95,59.5,-95</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>25.5 25</intersection>
<intersection>37 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37,-116.5,37,-95</points>
<intersection>-116.5 22</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>37,-116.5,44,-116.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>37 3</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>25.5,-96,25.5,-95</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-104,69.5,-104</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>65.5 3</intersection>
<intersection>69.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65.5,-126,65.5,-104</points>
<intersection>-126 4</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>65.5,-126,68,-126</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>69.5,-104,69.5,-104</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-104 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-254.5,69.5,-254.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>62 6</intersection>
<intersection>69.5 11</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>62,-267,62,-254.5</points>
<intersection>-267 9</intersection>
<intersection>-254.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>62,-267,71.5,-267</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>62 6</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>69.5,-255,69.5,-254.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-254.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-94,115.5,-94</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>115.5 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>115.5,-94.5,115.5,-94</points>
<connection>
<GID>49</GID>
<name>N_in0</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-101,69.5,-101</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>61 6</intersection>
<intersection>69.5 13</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>61,-128,61,-101</points>
<intersection>-128 9</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>61,-128,68,-128</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>61 6</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>69.5,-102,69.5,-101</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-101 1</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-103,98,-103</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>77 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>77,-115.5,77,-103</points>
<intersection>-115.5 6</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77,-115.5,95,-115.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>77 5</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-126.5,102.5,-126.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>74 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>74,-127,74,-126.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>-126.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-256,85.5,-251</points>
<intersection>-256 2</intersection>
<intersection>-251 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-251,95,-251</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection>
<intersection>89 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-256,85.5,-256</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>85.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>89,-259,89,-251</points>
<intersection>-259 6</intersection>
<intersection>-251 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89,-259,106,-259</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>89 5</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-104,121.5,-104</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>45</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-117.5,95,-117.5</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>92 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>92,-117.5,92,-105</points>
<intersection>-117.5 1</intersection>
<intersection>-105 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>92,-105,98,-105</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>92 4</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-124.5,101,-116.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>-124.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>101,-124.5,102.5,-124.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-125.5,121,-125.5</points>
<connection>
<GID>53</GID>
<name>N_in0</name></connection>
<connection>
<GID>48</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-25.5,166.5,-24</points>
<intersection>-25.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-24,166.5,-24</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-25.5,174.5,-25.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>166.5 0</intersection>
<intersection>168 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>168,-37.5,168,-25.5</points>
<intersection>-37.5 4</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>168,-37.5,169.5,-37.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>168 3</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-27.5,174.5,-27.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>156 9</intersection>
<intersection>170.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>170.5,-35.5,170.5,-27.5</points>
<intersection>-35.5 4</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>170.5,-35.5,176.5,-35.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>170.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>156,-29.5,156,-27.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173.5,-37.5,176.5,-37.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159,-50.5,177.5,-50.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>173.5 3</intersection>
<intersection>177.5 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>173.5,-58,173.5,-50.5</points>
<intersection>-58 4</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>173.5,-58,179.5,-58</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>173.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>177.5,-50.5,177.5,-50</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>176.5,-60,179.5,-60</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<connection>
<GID>68</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>180.5,-26.5,223.5,-26.5</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>74</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-60,169.5,-47.5</points>
<intersection>-60 4</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-47.5,177.5,-47.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection>
<intersection>177.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>169.5,-60,172.5,-60</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>177.5,-48,177.5,-47.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>-47.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-49,193.5,-44</points>
<intersection>-49 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-44,203,-44</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection>
<intersection>197 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-49,193.5,-49</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>193.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>197,-52,197,-44</points>
<intersection>-52 4</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>197,-52,207.5,-52</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>197 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-59.5,203,-59</points>
<intersection>-59.5 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-59.5,221.5,-59.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185.5,-59,203,-59</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>203 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>211.5,-52,214,-52</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209,-45,229,-45</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>77</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-54,153.5,-40.5</points>
<intersection>-54 1</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153.5,-54,214,-54</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>153.5 0</intersection>
<intersection>201 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153.5,-40.5,182.5,-40.5</points>
<intersection>153.5 0</intersection>
<intersection>182.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>182.5,-40.5,182.5,-36.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>-40.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>201,-54,201,-46</points>
<intersection>-54 1</intersection>
<intersection>-46 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>201,-46,203,-46</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>201 4</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221,-57.5,221,-53</points>
<intersection>-57.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221,-57.5,221.5,-57.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>221 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-53,221,-53</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>221 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-58.5,232.5,-58.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>78</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-88.5,170.5,-87</points>
<intersection>-88.5 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-87,170.5,-87</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170.5,-88.5,178.5,-88.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection>
<intersection>172 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>172,-100.5,172,-88.5</points>
<intersection>-100.5 6</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>172,-100.5,180.5,-100.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>172 5</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-90.5,178.5,-90.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>174.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>174.5,-98.5,174.5,-90.5</points>
<intersection>-98.5 4</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>174.5,-98.5,180.5,-98.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>174.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-113.5,181.5,-113.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>177.5 3</intersection>
<intersection>181.5 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>177.5,-121,177.5,-113.5</points>
<intersection>-121 4</intersection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>177.5,-121,183.5,-121</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>177.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>181.5,-113.5,181.5,-113</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>-113.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>184.5,-89.5,227.5,-89.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<connection>
<GID>102</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-110.5,181.5,-110.5</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>174 6</intersection>
<intersection>181.5 11</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>174,-123,174,-110.5</points>
<intersection>-123 9</intersection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>174,-123,183.5,-123</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>174 6</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>181.5,-111,181.5,-110.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-110.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-112,197.5,-107</points>
<intersection>-112 2</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197.5,-107,207,-107</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection>
<intersection>201 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-112,197.5,-112</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>197.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>201,-115,201,-107</points>
<intersection>-115 6</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>201,-115,218,-115</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>201 5</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-122.5,207,-122</points>
<intersection>-122.5 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-122.5,225.5,-122.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189.5,-122,207,-122</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-108,233,-108</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<connection>
<GID>105</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-117,157.5,-103.5</points>
<intersection>-117 1</intersection>
<intersection>-103.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-117,218,-117</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>157.5 0</intersection>
<intersection>205 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-103.5,186.5,-103.5</points>
<intersection>157.5 0</intersection>
<intersection>186.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>186.5,-103.5,186.5,-99.5</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>-103.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>205,-117,205,-109</points>
<intersection>-117 1</intersection>
<intersection>-109 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>205,-109,207,-109</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>205 4</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-120.5,225,-116</points>
<intersection>-120.5 1</intersection>
<intersection>-116 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-120.5,225.5,-120.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>224,-116,225,-116</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>231.5,-121.5,236.5,-121.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-266.5,95,-266</points>
<intersection>-266.5 1</intersection>
<intersection>-266 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-266.5,113.5,-266.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-266,95,-266</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-252,121,-252</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>44</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-261,45.5,-247.5</points>
<intersection>-261 1</intersection>
<intersection>-247.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-261,106,-261</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection>
<intersection>93 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-247.5,74.5,-247.5</points>
<intersection>45.5 0</intersection>
<intersection>74.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74.5,-247.5,74.5,-243.5</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>-247.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>93,-261,93,-253</points>
<intersection>-261 1</intersection>
<intersection>-253 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>93,-253,95,-253</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>93 4</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-264.5,113,-260</points>
<intersection>-264.5 1</intersection>
<intersection>-260 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,-264.5,113.5,-264.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112,-260,113,-260</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119.5,-265.5,124.5,-265.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>47</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>16.3888,171.387,156.24,25.2072</PageViewport>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>152.5,51.5</position>
<gparam>LABEL_TEXT green</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>288</ID>
<type>AA_LABEL</type>
<position>58,46</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>57.5,52</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>290</ID>
<type>AA_LABEL</type>
<position>56,70.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>56,59.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>56,34.5</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>57.5,23</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>140,67.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>299</ID>
<type>AA_LABEL</type>
<position>85,74.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>300</ID>
<type>AA_LABEL</type>
<position>84.5,67</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>301</ID>
<type>AA_LABEL</type>
<position>83.5,29</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>302</ID>
<type>AA_LABEL</type>
<position>83.5,21</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>304</ID>
<type>AA_LABEL</type>
<position>102.5,61</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>307</ID>
<type>AA_LABEL</type>
<position>148.5,69</position>
<gparam>LABEL_TEXT purple</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>15,-7</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>308</ID>
<type>AA_LABEL</type>
<position>101.5,50</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>42.5,-7.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>AA_LABEL</type>
<position>102,36</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>21.5,-7</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>145,28</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>48.5,-7</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>AA_LABEL</type>
<position>155.5,29.5</position>
<gparam>LABEL_TEXT brown</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_AND2</type>
<position>90,-15</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>97.5,-40</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>89.5,-69.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AE_OR2</type>
<position>103.5,-22.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND3</type>
<position>90,-28.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>66 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND3</type>
<position>89,-55</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>66 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_OR2</type>
<position>108,-62</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AO_XNOR2</type>
<position>67,-37.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AO_XNOR2</type>
<position>67,-43.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>121,-22.5</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>123,-40</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>GA_LED</type>
<position>127,-64.5</position>
<input>
<ID>N_in3</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_INVERTER</type>
<position>69,-31</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_INVERTER</type>
<position>73.5,-66.5</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_INVERTER</type>
<position>67.5,-51.5</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_INVERTER</type>
<position>69,-18.5</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>127.5,-21.5</position>
<gparam>LABEL_TEXT A>B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>129.5,-39</position>
<gparam>LABEL_TEXT A=B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>133,-63.5</position>
<gparam>LABEL_TEXT AB</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_TOGGLE</type>
<position>15.5,-10</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_TOGGLE</type>
<position>21,-10</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_TOGGLE</type>
<position>43,-10.5</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_TOGGLE</type>
<position>48.5,-10.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>49,52.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>49,46</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>17.5,93</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>35.5,92</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>23.5,92.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>41,92</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_AND2</type>
<position>85,74</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>102,49</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND2</type>
<position>84,20.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_OR2</type>
<position>140.5,67</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_OR2</type>
<position>145,27.5</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>158,67</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>GA_LED</type>
<position>160,49.5</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>164,25</position>
<input>
<ID>N_in3</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_INVERTER</type>
<position>57,59</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_INVERTER</type>
<position>58.5,23</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_INVERTER</type>
<position>57,34</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_INVERTER</type>
<position>56.5,70</position>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>164.5,68</position>
<gparam>LABEL_TEXT A>B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>166.5,50.5</position>
<gparam>LABEL_TEXT A=B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>170,26</position>
<gparam>LABEL_TEXT AB</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_TOGGLE</type>
<position>18,88</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_TOGGLE</type>
<position>23.5,87.5</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_TOGGLE</type>
<position>35,87.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_TOGGLE</type>
<position>40.5,87.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>182</ID>
<type>AI_XOR2</type>
<position>49,52</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_INVERTER</type>
<position>58.5,51.5</position>
<input>
<ID>IN_0</ID>96 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>186</ID>
<type>AI_XOR2</type>
<position>49,45.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_INVERTER</type>
<position>59,45.5</position>
<input>
<ID>IN_0</ID>97 </input>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>84.5,66</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_AND2</type>
<position>103,60.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND2</type>
<position>84,28.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_AND2</type>
<position>102.5,36</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>15</ID>
<points>48.5,-55,48.5,-12.5</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>-55 30</intersection>
<intersection>-42.5 28</intersection>
<intersection>-31 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>48.5,-31,66,-31</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>48.5 15</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>48.5,-42.5,64,-42.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>48.5 15</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>48.5,-55,86,-55</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>48.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>15</ID>
<points>43.5,-70.5,43.5,-12.5</points>
<intersection>-70.5 32</intersection>
<intersection>-38.5 30</intersection>
<intersection>-18.5 28</intersection>
<intersection>-12.5 33</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>43.5,-18.5,66,-18.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>43.5 15</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>43.5,-38.5,64,-38.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>43.5 15</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>43.5,-70.5,86.5,-70.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>43.5 15</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>43,-12.5,43.5,-12.5</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>43.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-51.5,20,-26.5</points>
<intersection>-51.5 11</intersection>
<intersection>-44.5 13</intersection>
<intersection>-26.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>20,-26.5,87,-26.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection>
<intersection>21 14</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>20,-51.5,64.5,-51.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>20,-44.5,64,-44.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>21,-26.5,21,-12</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-66.5,16.5,-12</points>
<intersection>-66.5 13</intersection>
<intersection>-36.5 11</intersection>
<intersection>-14 9</intersection>
<intersection>-12 14</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>16.5,-14,87,-14</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>16.5,-36.5,64,-36.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>16.5,-66.5,70.5,-66.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>15.5,-12,16.5,-12</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-21.5,96.5,-15</points>
<intersection>-21.5 1</intersection>
<intersection>-15 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-21.5,100.5,-21.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>93,-15,96.5,-15</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>99.5,-61,99.5,-55</points>
<intersection>-61 4</intersection>
<intersection>-55 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>99.5,-61,105,-61</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>99.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>92,-55,99.5,-55</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>99.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-69.5,99.5,-63</points>
<intersection>-69.5 4</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-63,105,-63</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>92.5,-69.5,99.5,-69.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-41,94.5,-41</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>85 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85,-43.5,85,-41</points>
<intersection>-43.5 4</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>70,-43.5,85,-43.5</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>85 3</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-23.5,100.5,-23.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>96.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>96.5,-28.5,96.5,-23.5</points>
<intersection>-28.5 8</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>93,-28.5,96.5,-28.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>96.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-57,83.5,-30.5</points>
<intersection>-57 5</intersection>
<intersection>-37.5 2</intersection>
<intersection>-37 6</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-30.5,87,-30.5</points>
<connection>
<GID>123</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-37.5,83.5,-37.5</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>83.5,-57,86,-57</points>
<connection>
<GID>124</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>83.5,-37,94.5,-37</points>
<intersection>83.5 0</intersection>
<intersection>94.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>94.5,-39,94.5,-37</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-37 6</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-22.5,120,-22.5</points>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<connection>
<GID>122</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-62,127,-62</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>127 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>127,-63.5,127,-62</points>
<connection>
<GID>130</GID>
<name>N_in3</name></connection>
<intersection>-62 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-40,122,-40</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-18.5,87,-18.5</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>87 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>87,-18.5,87,-16</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-68.5,80.5,-66.5</points>
<intersection>-68.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-68.5,86.5,-68.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-66.5,80.5,-66.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-31,79.5,-28.5</points>
<intersection>-31 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-28.5,87,-28.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-31,79.5,-31</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-53,78,-51.5</points>
<intersection>-53 1</intersection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-53,86,-53</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-51.5,78,-51.5</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>15</ID>
<points>40.5,27.5,40.5,85.5</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>27.5 30</intersection>
<intersection>44.5 32</intersection>
<intersection>59 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>40.5,59,54,59</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>40.5 15</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>40.5,27.5,81,27.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>40.5 15</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>40.5,44.5,46,44.5</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>40.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>15</ID>
<points>35,20,35,85.5</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>20 32</intersection>
<intersection>51 35</intersection>
<intersection>70 28</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>35,70,53.5,70</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>35 15</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>35,20,81,20</points>
<intersection>35 15</intersection>
<intersection>81 37</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>35,51,46,51</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>35 15</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>81,19.5,81,20</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>20 32</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,34,23.5,85.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>34 11</intersection>
<intersection>46.5 17</intersection>
<intersection>67 19</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>23.5,34,54,34</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>23.5,46.5,46,46.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>23.5,67,81.5,67</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,23,18,86</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>23 13</intersection>
<intersection>53 17</intersection>
<intersection>75 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>18,75,82,75</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>18,23,55.5,23</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>18,53,46,53</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,68,98,74</points>
<intersection>68 1</intersection>
<intersection>74 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,68,137.5,68</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>88,74,98,74</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>108,28.5,108,36</points>
<intersection>28.5 4</intersection>
<intersection>36 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>108,28.5,142,28.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>108 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>105.5,36,108,36</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>108 3</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,20.5,101,26.5</points>
<intersection>20.5 4</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,26.5,142,26.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>87,20.5,101,20.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122,66,137.5,66</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>122 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>122,60.5,122,66</points>
<intersection>60.5 12</intersection>
<intersection>66 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>106,60.5,122,60.5</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>122 9</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,35,89.5,59.5</points>
<intersection>35 16</intersection>
<intersection>50 6</intersection>
<intersection>52.5 13</intersection>
<intersection>59.5 15</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,50,99,50</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>61.5,52.5,89.5,52.5</points>
<intersection>61.5 17</intersection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>89.5,59.5,100,59.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>89.5,35,99.5,35</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>61.5,51.5,61.5,52.5</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>52.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>143.5,67,157,67</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<connection>
<GID>167</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148,27.5,164,27.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>164 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>164,26,164,27.5</points>
<connection>
<GID>169</GID>
<name>N_in3</name></connection>
<intersection>27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,49,159,49</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>159 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>159,49,159,49.5</points>
<connection>
<GID>168</GID>
<name>N_in0</name></connection>
<intersection>49 1</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,70,60.5,70</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>60.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>60.5,70,60.5,73</points>
<intersection>70 1</intersection>
<intersection>73 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>60.5,73,82,73</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>60.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,21.5,64,23</points>
<intersection>21.5 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,21.5,81,21.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,23,64,23</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,59,73.5,65</points>
<intersection>59 4</intersection>
<intersection>65 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>73.5,65,81.5,65</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>60,59,73.5,59</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,29.5,63.5,34</points>
<intersection>29.5 4</intersection>
<intersection>34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,34,63.5,34</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>63.5,29.5,81,29.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,51.5,55.5,51.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>52 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>52,51.5,52,52</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,45.5,56,45.5</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,45.5,88,48</points>
<intersection>45.5 2</intersection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,48,99,48</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62,45.5,88,45.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,66,100,66</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>100 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>100,61.5,100,66</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>66 1</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,37,99.5,37</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>87 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>87,28.5,87,37</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>37 1</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>-86.4408,45.5399,-34.0556,-9.21574</PageViewport>
<gate>
<ID>193</ID>
<type>GA_LED</type>
<position>18.5,4</position>
<input>
<ID>N_in0</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>29.5,8</position>
<gparam>LABEL_TEXT AND</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-35.5,29.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>195</ID>
<type>GA_LED</type>
<position>18.5,-4</position>
<input>
<ID>N_in1</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>GA_LED</type>
<position>18.5,-9</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AE_OR2</type>
<position>10.5,-4</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-32.5,29.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>198</ID>
<type>AE_OR2</type>
<position>10.5,-9</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AI_XOR2</type>
<position>10.5,-17</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-26.5,29.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>GA_LED</type>
<position>18.5,-17</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>GA_LED</type>
<position>18.5,-22</position>
<input>
<ID>N_in0</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AI_XOR2</type>
<position>10.5,-22</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>29.5,-5</position>
<gparam>LABEL_TEXT OR</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>AA_LABEL</type>
<position>29.5,-18</position>
<gparam>LABEL_TEXT XOR</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>-23.5,29.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>-23.5,32</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>-26.5,32</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_LABEL</type>
<position>-32.5,32</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_LABEL</type>
<position>-35.5,32</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>9.5,9.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND2</type>
<position>10.5,4</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>GA_LED</type>
<position>18.5,9</position>
<input>
<ID>N_in0</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-16,-23.5,27.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-16 7</intersection>
<intersection>-3 5</intersection>
<intersection>10.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-23.5,10.5,6.5,10.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-23.5,-3,7.5,-3</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-23.5,-16,7.5,-16</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-21,-26.5,27.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-21 7</intersection>
<intersection>-8 5</intersection>
<intersection>5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-26.5,5,7.5,5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-26.5,-8,7.5,-8</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-26.5,-21,7.5,-21</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-18,-32.5,27.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-18 7</intersection>
<intersection>-5 5</intersection>
<intersection>8.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-32.5,8.5,6.5,8.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-32.5,-5,7.5,-5</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-32.5,-18,7.5,-18</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-23,-35.5,27.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-23 7</intersection>
<intersection>-10 5</intersection>
<intersection>3 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-35.5,3,7.5,3</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-35.5,-10,7.5,-10</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-35.5,-23,7.5,-23</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,9.5,17.5,9.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>17.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>17.5,9,17.5,9.5</points>
<connection>
<GID>192</GID>
<name>N_in0</name></connection>
<intersection>9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,4,17.5,4</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<connection>
<GID>193</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-4,19.5,-4</points>
<connection>
<GID>197</GID>
<name>OUT</name></connection>
<connection>
<GID>195</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-9,17.5,-9</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<connection>
<GID>196</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-17,17.5,-17</points>
<connection>
<GID>200</GID>
<name>N_in0</name></connection>
<connection>
<GID>199</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-22,17.5,-22</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<connection>
<GID>201</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-406.472,139.845,-116.099,-163.668</PageViewport>
<gate>
<ID>388</ID>
<type>AA_INVERTER</type>
<position>0,-177</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>389</ID>
<type>AA_INVERTER</type>
<position>1.5,-213</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>390</ID>
<type>AA_INVERTER</type>
<position>0,-202</position>
<input>
<ID>IN_0</ID>118 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>391</ID>
<type>AA_INVERTER</type>
<position>-0.5,-166</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>399</ID>
<type>AI_XOR2</type>
<position>-8,-184</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>AA_INVERTER</type>
<position>1.5,-184.5</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>401</ID>
<type>AI_XOR2</type>
<position>-8,-190.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>AA_INVERTER</type>
<position>2,-190.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>403</ID>
<type>AA_AND2</type>
<position>27.5,-170</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_AND2</type>
<position>46,-175.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>27,-207.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>45.5,-200</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_LABEL</type>
<position>33,-146.5</position>
<gparam>LABEL_TEXT 2 bit Comaparator</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>409</ID>
<type>AE_MUX_4x1</type>
<position>120.5,-119</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>153 </input>
<output>
<ID>OUT</ID>168 </output>
<input>
<ID>SEL_0</ID>165 </input>
<input>
<ID>SEL_1</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>411</ID>
<type>AI_MUX_8x1</type>
<position>120.5,-89</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>175 </input>
<input>
<ID>IN_2</ID>178 </input>
<input>
<ID>IN_3</ID>184 </input>
<input>
<ID>IN_4</ID>185 </input>
<input>
<ID>IN_5</ID>186 </input>
<output>
<ID>OUT</ID>170 </output>
<input>
<ID>SEL_0</ID>165 </input>
<input>
<ID>SEL_1</ID>166 </input>
<input>
<ID>SEL_2</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>413</ID>
<type>AI_MUX_8x1</type>
<position>120.5,-73</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>174 </input>
<input>
<ID>IN_2</ID>177 </input>
<input>
<ID>IN_3</ID>179 </input>
<input>
<ID>IN_4</ID>181 </input>
<input>
<ID>IN_5</ID>180 </input>
<output>
<ID>OUT</ID>171 </output>
<input>
<ID>SEL_0</ID>165 </input>
<input>
<ID>SEL_1</ID>166 </input>
<input>
<ID>SEL_2</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>415</ID>
<type>GA_LED</type>
<position>-30,-7</position>
<input>
<ID>N_in3</ID>168 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>416</ID>
<type>GA_LED</type>
<position>-23,-7</position>
<input>
<ID>N_in3</ID>170 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>417</ID>
<type>GA_LED</type>
<position>-16,-7</position>
<input>
<ID>N_in3</ID>171 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>418</ID>
<type>AA_LABEL</type>
<position>-30.5,-9</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>419</ID>
<type>AA_LABEL</type>
<position>-23.5,-9</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>420</ID>
<type>AA_LABEL</type>
<position>-16,-9</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>421</ID>
<type>AA_LABEL</type>
<position>-16,-11</position>
<gparam>LABEL_TEXT A>B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>AA_LABEL</type>
<position>-30.5,-11</position>
<gparam>LABEL_TEXT AB</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>AA_LABEL</type>
<position>-23.5,-11</position>
<gparam>LABEL_TEXT A=B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>425</ID>
<type>AA_AND2</type>
<position>102,-73.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>427</ID>
<type>AE_OR2</type>
<position>102,-69</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>AI_XOR2</type>
<position>102.5,-64.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>AA_AND2</type>
<position>101.5,-96.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>431</ID>
<type>AE_OR2</type>
<position>101.5,-92</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>432</ID>
<type>AI_XOR2</type>
<position>102,-87.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>261</ID>
<type>AI_XOR2</type>
<position>32,-49</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_AND2</type>
<position>25.5,-60.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_SMALL_INVERTER</type>
<position>17.5,-61.5</position>
<input>
<ID>IN_0</ID>118 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>264</ID>
<type>AI_XOR2</type>
<position>26.5,-73</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>28.5,-83</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>AE_SMALL_INVERTER</type>
<position>20.5,-84</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>267</ID>
<type>AI_XOR2</type>
<position>52,-69</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>63,-77</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_SMALL_INVERTER</type>
<position>55.5,-76</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_OR2</type>
<position>70.5,-83</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>17,-60.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>AA_LABEL</type>
<position>20.5,-83.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>AA_LABEL</type>
<position>55,-75.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>279</ID>
<type>AA_LABEL</type>
<position>32,-48.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>280</ID>
<type>AA_LABEL</type>
<position>32,-37.5</position>
<gparam>LABEL_TEXT 2 bit Substraction</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>AA_LABEL</type>
<position>13.5,-42.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>282</ID>
<type>AA_LABEL</type>
<position>16.5,-48.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>AA_LABEL</type>
<position>16,-68.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>AA_LABEL</type>
<position>21,-72.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>AA_LABEL</type>
<position>26.5,-72.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_LABEL</type>
<position>52,-68.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>297</ID>
<type>AA_LABEL</type>
<position>25.5,-60</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>298</ID>
<type>AA_LABEL</type>
<position>28,-82.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>303</ID>
<type>AA_LABEL</type>
<position>62.5,-76.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>305</ID>
<type>AA_LABEL</type>
<position>70.5,-82.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>313</ID>
<type>AI_XOR2</type>
<position>24,-103</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_AND2</type>
<position>8.5,-126.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AI_XOR2</type>
<position>34,-112</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>32.5,-136</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>AI_XOR2</type>
<position>62.5,-113</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>140 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_AND2</type>
<position>59.5,-125.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>140 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_OR2</type>
<position>67,-134.5</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_LABEL</type>
<position>33.5,-94.5</position>
<gparam>LABEL_TEXT 2 bit Addition</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>333</ID>
<type>AA_LABEL</type>
<position>24,-102.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>334</ID>
<type>AA_LABEL</type>
<position>34,-111.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>335</ID>
<type>AA_LABEL</type>
<position>8,-126</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>336</ID>
<type>AA_LABEL</type>
<position>59.5,-125</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>337</ID>
<type>AA_LABEL</type>
<position>62.5,-112.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>338</ID>
<type>AA_LABEL</type>
<position>32.5,-135.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>339</ID>
<type>AA_LABEL</type>
<position>67,-134</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>341</ID>
<type>AA_TOGGLE</type>
<position>-32.5,-22</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>342</ID>
<type>AA_TOGGLE</type>
<position>-29,-22</position>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_TOGGLE</type>
<position>-24,-22</position>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_TOGGLE</type>
<position>-21,-22</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_TOGGLE</type>
<position>-16,-22</position>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>346</ID>
<type>AA_TOGGLE</type>
<position>-13,-22</position>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>347</ID>
<type>AA_TOGGLE</type>
<position>-10,-22</position>
<output>
<ID>OUT_0</ID>165 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_LABEL</type>
<position>-32.5,-19.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>AA_LABEL</type>
<position>-28.5,-19.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>AA_LABEL</type>
<position>-24.5,-19.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>AA_LABEL</type>
<position>-20.5,-19.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>353</ID>
<type>AA_LABEL</type>
<position>-13,-19.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>AA_LABEL</type>
<position>-9.5,-19.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>AA_LABEL</type>
<position>-16,-19.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>357</ID>
<type>AA_LABEL</type>
<position>1,-190</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>358</ID>
<type>AA_LABEL</type>
<position>0.5,-184</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>359</ID>
<type>AA_LABEL</type>
<position>-1,-165.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>360</ID>
<type>AA_LABEL</type>
<position>-1,-176.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>361</ID>
<type>AA_LABEL</type>
<position>-1,-201.5</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>0.5,-213</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>363</ID>
<type>AA_LABEL</type>
<position>83,-168.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_LABEL</type>
<position>28,-161.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>27.5,-169</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>366</ID>
<type>AA_LABEL</type>
<position>26.5,-207</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>367</ID>
<type>AA_LABEL</type>
<position>26.5,-215</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>368</ID>
<type>AA_LABEL</type>
<position>45.5,-175</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>370</ID>
<type>AA_LABEL</type>
<position>44.5,-186</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>371</ID>
<type>AA_LABEL</type>
<position>45,-200</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>372</ID>
<type>AA_LABEL</type>
<position>88,-208</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>374</ID>
<type>AA_LABEL</type>
<position>-8,-183.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>375</ID>
<type>AA_LABEL</type>
<position>-8,-190</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>380</ID>
<type>AA_AND2</type>
<position>28,-162</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>AA_AND2</type>
<position>45,-187</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_AND2</type>
<position>27,-215.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>AE_OR2</type>
<position>83.5,-169</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>AE_OR2</type>
<position>88,-208.5</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29,-44,94,-44</points>
<intersection>-29 3</intersection>
<intersection>27.5 11</intersection>
<intersection>94 25</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-29,-202,-29,-24</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>-202 22</intersection>
<intersection>-189.5 20</intersection>
<intersection>-169 18</intersection>
<intersection>-127.5 16</intersection>
<intersection>-102 14</intersection>
<intersection>-61.5 4</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-29,-61.5,15.5,-61.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>-29 3</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>27.5,-48,27.5,-44</points>
<intersection>-48 24</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-29,-102,21,-102</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>-29 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-29,-127.5,5.5,-127.5</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>-29 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-29,-169,24.5,-169</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>-29 3</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-29,-189.5,-11,-189.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>-29 3</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-29,-202,-3,-202</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-29 3</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>27.5,-48,29,-48</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>27.5 11</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>94,-72.5,94,-44</points>
<intersection>-72.5 30</intersection>
<intersection>-68 28</intersection>
<intersection>-63.5 26</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>94,-63.5,99.5,-63.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>94 25</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>94,-68,99,-68</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>94 25</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>94,-72.5,99,-72.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>94 25</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-54.5,95,-54.5</points>
<intersection>-21 3</intersection>
<intersection>95 24</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-21,-208.5,-21,-24</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>-208.5 23</intersection>
<intersection>-191.5 21</intersection>
<intersection>-177 19</intersection>
<intersection>-125.5 17</intersection>
<intersection>-104 15</intersection>
<intersection>-59.5 4</intersection>
<intersection>-54.5 1</intersection>
<intersection>-50 26</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-21,-59.5,22.5,-59.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-21 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-21,-104,21,-104</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>-21 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-21,-125.5,5.5,-125.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>-21 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-21,-177,-3,-177</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-21 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-21,-191.5,-11,-191.5</points>
<connection>
<GID>401</GID>
<name>IN_1</name></connection>
<intersection>-21 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-21,-208.5,24,-208.5</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>-21 3</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>95,-74.5,95,-54.5</points>
<intersection>-74.5 32</intersection>
<intersection>-70 30</intersection>
<intersection>-65.5 27</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>-21,-50,29,-50</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>-21 3</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>95,-65.5,99.5,-65.5</points>
<connection>
<GID>429</GID>
<name>IN_1</name></connection>
<intersection>95 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>95,-70,99,-70</points>
<connection>
<GID>427</GID>
<name>IN_1</name></connection>
<intersection>95 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>95,-74.5,99,-74.5</points>
<connection>
<GID>425</GID>
<name>IN_1</name></connection>
<intersection>95 24</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-61.5,22.5,-61.5</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<connection>
<GID>262</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-24,-74,23.5,-74</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>-24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-24,-216.5,-24,-24</points>
<connection>
<GID>343</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 18</intersection>
<intersection>-185 16</intersection>
<intersection>-166 14</intersection>
<intersection>-135 12</intersection>
<intersection>-113 10</intersection>
<intersection>-88.5 20</intersection>
<intersection>-82 4</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-24,-82,25.5,-82</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-24 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-24,-113,31,-113</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>-24 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-24,-135,29.5,-135</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>-24 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-24,-166,-3.5,-166</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>-24 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-24,-185,-11,-185</points>
<connection>
<GID>399</GID>
<name>IN_1</name></connection>
<intersection>-24 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-24,-216.5,24,-216.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>-24 3</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-24,-88.5,99,-88.5</points>
<connection>
<GID>432</GID>
<name>IN_1</name></connection>
<intersection>-24 3</intersection>
<intersection>93 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>93,-97.5,93,-88.5</points>
<intersection>-97.5 25</intersection>
<intersection>-93 22</intersection>
<intersection>-88.5 20</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>93,-93,98.5,-93</points>
<connection>
<GID>431</GID>
<name>IN_1</name></connection>
<intersection>93 21</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>93,-97.5,98.5,-97.5</points>
<connection>
<GID>430</GID>
<name>IN_1</name></connection>
<intersection>93 21</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-84,25.5,-84</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<connection>
<GID>265</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-49,109,-49</points>
<connection>
<GID>261</GID>
<name>OUT</name></connection>
<intersection>109 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>109,-76.5,109,-49</points>
<intersection>-76.5 9</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>109,-76.5,117.5,-76.5</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>109 8</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-213,-32.5,-24</points>
<connection>
<GID>341</GID>
<name>OUT_0</name></connection>
<intersection>-213 19</intersection>
<intersection>-183 17</intersection>
<intersection>-161 15</intersection>
<intersection>-137 13</intersection>
<intersection>-111 22</intersection>
<intersection>-86.5 11</intersection>
<intersection>-84 4</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-70.5,23.5,-70.5</points>
<intersection>-32.5 0</intersection>
<intersection>23.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-32.5,-84,18.5,-84</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>23.5,-72,23.5,-70.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-32.5,-86.5,99,-86.5</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection>
<intersection>92 23</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-32.5,-137,29.5,-137</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-32.5,-161,25,-161</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-32.5,-183,-11,-183</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-32.5,-213,-1.5,-213</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-32.5,-111,31,-111</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>92,-95.5,92,-86.5</points>
<intersection>-95.5 26</intersection>
<intersection>-91 24</intersection>
<intersection>-86.5 11</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>92,-91,98.5,-91</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>92 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>92,-95.5,98.5,-95.5</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>92 23</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-73,39.5,-68</points>
<intersection>-73 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-68,49,-68</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection>
<intersection>43 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-73,39.5,-73</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43,-76,43,-68</points>
<intersection>-76 4</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43,-76,53.5,-76</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>43 3</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-84,49,-83</points>
<intersection>-84 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-84,67.5,-84</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-83,49,-83</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-76,60,-76</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<connection>
<GID>268</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-78,-0.5,-64.5</points>
<intersection>-78 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-78,60,-78</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>-0.5 0</intersection>
<intersection>47 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-64.5,28.5,-64.5</points>
<intersection>-0.5 0</intersection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28.5,-64.5,28.5,-60.5</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-64.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>47,-78,47,-70</points>
<intersection>-78 1</intersection>
<intersection>-70 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>47,-70,49,-70</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<intersection>47 4</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-82,67,-77</points>
<intersection>-82 1</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-82,67.5,-82</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,-77,67,-77</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-112,59.5,-112</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>38.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>38.5,-124.5,38.5,-112</points>
<intersection>-124.5 6</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>38.5,-124.5,56.5,-124.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>38.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-135.5,64,-135.5</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>35.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>35.5,-136,35.5,-135.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>-135.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-126.5,56.5,-126.5</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-126.5,53.5,-114</points>
<intersection>-126.5 1</intersection>
<intersection>-114 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>53.5,-114,59.5,-114</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>53.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-133.5,62.5,-125.5</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<intersection>-133.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>62.5,-133.5,64,-133.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-168,41,-162</points>
<intersection>-168 1</intersection>
<intersection>-162 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-168,80.5,-168</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>31,-162,41,-162</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>51,-207.5,51,-200</points>
<intersection>-207.5 4</intersection>
<intersection>-200 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51,-207.5,85,-207.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>51 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>48.5,-200,51,-200</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<intersection>51 3</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-215.5,44,-209.5</points>
<intersection>-215.5 4</intersection>
<intersection>-209.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-209.5,85,-209.5</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>30,-215.5,44,-215.5</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-170,80.5,-170</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>65 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>65,-175.5,65,-170</points>
<intersection>-175.5 12</intersection>
<intersection>-170 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>49,-175.5,65,-175.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>65 9</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-201,32.5,-176.5</points>
<intersection>-201 16</intersection>
<intersection>-186 6</intersection>
<intersection>-183.5 13</intersection>
<intersection>-176.5 15</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>32.5,-186,42,-186</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>4.5,-183.5,32.5,-183.5</points>
<intersection>4.5 17</intersection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>32.5,-176.5,43,-176.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>32.5,-201,42.5,-201</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>4.5,-184.5,4.5,-183.5</points>
<connection>
<GID>400</GID>
<name>OUT_0</name></connection>
<intersection>-183.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91,-208.5,117.5,-208.5</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<intersection>117.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>117.5,-208.5,117.5,-118</points>
<connection>
<GID>409</GID>
<name>IN_2</name></connection>
<intersection>-208.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-166,3.5,-166</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<intersection>3.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>3.5,-166,3.5,-163</points>
<intersection>-166 1</intersection>
<intersection>-163 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>3.5,-163,25,-163</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>3.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-214.5,7,-213</points>
<intersection>-214.5 1</intersection>
<intersection>-213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-214.5,24,-214.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-213,7,-213</points>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-177,16.5,-171</points>
<intersection>-177 4</intersection>
<intersection>-171 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>16.5,-171,24.5,-171</points>
<connection>
<GID>403</GID>
<name>IN_1</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>3,-177,16.5,-177</points>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-206.5,6.5,-202</points>
<intersection>-206.5 4</intersection>
<intersection>-202 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>3,-202,6.5,-202</points>
<connection>
<GID>390</GID>
<name>OUT_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>6.5,-206.5,24,-206.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,-184.5,-1.5,-184.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>-5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-5,-184.5,-5,-184</points>
<connection>
<GID>399</GID>
<name>OUT</name></connection>
<intersection>-184.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,-190.5,-1,-190.5</points>
<connection>
<GID>401</GID>
<name>OUT</name></connection>
<connection>
<GID>402</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-190.5,31,-188</points>
<intersection>-190.5 2</intersection>
<intersection>-188 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-188,42,-188</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-190.5,31,-190.5</points>
<connection>
<GID>402</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-170,43,-170</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<intersection>43 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43,-174.5,43,-170</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-170 1</intersection></vsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-199,42.5,-199</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>30 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>30,-207.5,30,-199</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>-199 1</intersection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-114,121.5,-28</points>
<connection>
<GID>409</GID>
<name>SEL_0</name></connection>
<connection>
<GID>411</GID>
<name>SEL_0</name></connection>
<connection>
<GID>413</GID>
<name>SEL_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-10,-28,-10,-24</points>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-10,-28,121.5,-28</points>
<intersection>-10 1</intersection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-114,120.5,-30.5</points>
<connection>
<GID>409</GID>
<name>SEL_1</name></connection>
<connection>
<GID>411</GID>
<name>SEL_1</name></connection>
<connection>
<GID>413</GID>
<name>SEL_1</name></connection>
<intersection>-30.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-13,-30.5,-13,-24</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13,-30.5,120.5,-30.5</points>
<intersection>-13 1</intersection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-83.5,119.5,-32.5</points>
<connection>
<GID>411</GID>
<name>SEL_2</name></connection>
<connection>
<GID>413</GID>
<name>SEL_2</name></connection>
<intersection>-32.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-16,-32.5,-16,-24</points>
<connection>
<GID>345</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-16,-32.5,119.5,-32.5</points>
<intersection>-16 1</intersection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-6,-30,11.5</points>
<connection>
<GID>415</GID>
<name>N_in3</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,11.5,141,11.5</points>
<intersection>-30 0</intersection>
<intersection>141 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>141,-119,141,11.5</points>
<intersection>-119 3</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123.5,-119,141,-119</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<intersection>141 2</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23,1,138.5,1</points>
<intersection>-23 3</intersection>
<intersection>138.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-23,-6,-23,1</points>
<connection>
<GID>416</GID>
<name>N_in3</name></connection>
<intersection>1 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>138.5,-89,138.5,1</points>
<intersection>-89 5</intersection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>123.5,-89,138.5,-89</points>
<connection>
<GID>411</GID>
<name>OUT</name></connection>
<intersection>138.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,-2.5,132.5,-2.5</points>
<intersection>-16 7</intersection>
<intersection>132.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132.5,-73,132.5,-2.5</points>
<intersection>-73 4</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>123.5,-73,132.5,-73</points>
<connection>
<GID>413</GID>
<name>OUT</name></connection>
<intersection>132.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-16,-6,-16,-2.5</points>
<connection>
<GID>417</GID>
<name>N_in3</name></connection>
<intersection>-2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-92.5,108,-68.5</points>
<intersection>-92.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-68.5,108,-68.5</points>
<intersection>55 3</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,-92.5,117.5,-92.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,-69,55,-68.5</points>
<connection>
<GID>267</GID>
<name>OUT</name></connection>
<intersection>-68.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-122,101,-83</points>
<intersection>-122 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-83,101,-83</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-122,117.5,-122</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-103,109.5,-75.5</points>
<intersection>-103 1</intersection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-103,109.5,-103</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-75.5,117.5,-75.5</points>
<connection>
<GID>413</GID>
<name>IN_1</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-113,110.5,-91.5</points>
<intersection>-113 2</intersection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-91.5,117.5,-91.5</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-113,110.5,-113</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-134.5,110.5,-120</points>
<intersection>-134.5 2</intersection>
<intersection>-120 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-120,117.5,-120</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-134.5,110.5,-134.5</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-169,110.5,-74.5</points>
<intersection>-169 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-169,110.5,-169</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-74.5,117.5,-74.5</points>
<connection>
<GID>413</GID>
<name>IN_2</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-187,107,-91</points>
<intersection>-187 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-91,117.5,-91</points>
<intersection>107 0</intersection>
<intersection>117.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-187,107,-187</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117.5,-91,117.5,-90.5</points>
<connection>
<GID>411</GID>
<name>IN_2</name></connection>
<intersection>-91 1</intersection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-73.5,117.5,-73.5</points>
<connection>
<GID>413</GID>
<name>IN_3</name></connection>
<connection>
<GID>425</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-71.5,111.5,-64.5</points>
<intersection>-71.5 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-71.5,117.5,-71.5</points>
<connection>
<GID>413</GID>
<name>IN_5</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-64.5,111.5,-64.5</points>
<connection>
<GID>429</GID>
<name>OUT</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-72.5,111,-69</points>
<intersection>-72.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-72.5,117.5,-72.5</points>
<connection>
<GID>413</GID>
<name>IN_4</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,-69,111,-69</points>
<connection>
<GID>427</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-96.5,112,-89.5</points>
<intersection>-96.5 2</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-89.5,117.5,-89.5</points>
<connection>
<GID>411</GID>
<name>IN_3</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-96.5,112,-96.5</points>
<connection>
<GID>430</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-88.5,117.5,-88.5</points>
<connection>
<GID>411</GID>
<name>IN_4</name></connection>
<intersection>106.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>106.5,-92,106.5,-88.5</points>
<intersection>-92 4</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-92,106.5,-92</points>
<connection>
<GID>431</GID>
<name>OUT</name></connection>
<intersection>106.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-87.5,117.5,-87.5</points>
<connection>
<GID>411</GID>
<name>IN_5</name></connection>
<connection>
<GID>432</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-191.385,206.615,-16.9642,24.3026</PageViewport>
<gate>
<ID>433</ID>
<type>AA_INVERTER</type>
<position>44,-48</position>
<input>
<ID>IN_0</ID>188 </input>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>434</ID>
<type>AA_INVERTER</type>
<position>45.5,-84</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>435</ID>
<type>AA_INVERTER</type>
<position>44,-73</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>212 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>436</ID>
<type>AA_INVERTER</type>
<position>41,-37</position>
<input>
<ID>IN_0</ID>190 </input>
<output>
<ID>OUT_0</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>437</ID>
<type>AI_XOR2</type>
<position>36,-55</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>438</ID>
<type>AA_INVERTER</type>
<position>45.5,-55.5</position>
<input>
<ID>IN_0</ID>213 </input>
<output>
<ID>OUT_0</ID>207 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>439</ID>
<type>AI_XOR2</type>
<position>36,-61.5</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_INVERTER</type>
<position>46,-61.5</position>
<input>
<ID>IN_0</ID>214 </input>
<output>
<ID>OUT_0</ID>215 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>441</ID>
<type>AA_AND2</type>
<position>71.5,-41</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>442</ID>
<type>AA_AND2</type>
<position>90,-46.5</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>AA_AND2</type>
<position>71,-78.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>444</ID>
<type>AA_AND2</type>
<position>89.5,-71</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_LABEL</type>
<position>77,-17.5</position>
<gparam>LABEL_TEXT 2 bit Comaparator</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>446</ID>
<type>AE_MUX_4x1</type>
<position>164.5,10</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>228 </input>
<input>
<ID>IN_2</ID>208 </input>
<input>
<ID>IN_3</ID>237 </input>
<output>
<ID>OUT</ID>221 </output>
<input>
<ID>SEL_0</ID>218 </input>
<input>
<ID>SEL_1</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>447</ID>
<type>AI_MUX_8x1</type>
<position>164.5,40</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>227 </input>
<input>
<ID>IN_2</ID>230 </input>
<input>
<ID>IN_3</ID>234 </input>
<input>
<ID>IN_4</ID>243 </input>
<input>
<ID>IN_5</ID>242 </input>
<input>
<ID>IN_6</ID>238 </input>
<input>
<ID>IN_7</ID>238 </input>
<output>
<ID>OUT</ID>222 </output>
<input>
<ID>SEL_0</ID>218 </input>
<input>
<ID>SEL_1</ID>219 </input>
<input>
<ID>SEL_2</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>448</ID>
<type>AI_MUX_8x1</type>
<position>164.5,56</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>226 </input>
<input>
<ID>IN_2</ID>229 </input>
<input>
<ID>IN_3</ID>231 </input>
<input>
<ID>IN_4</ID>241 </input>
<input>
<ID>IN_5</ID>240 </input>
<input>
<ID>IN_6</ID>239 </input>
<input>
<ID>IN_7</ID>239 </input>
<output>
<ID>OUT</ID>223 </output>
<input>
<ID>SEL_0</ID>218 </input>
<input>
<ID>SEL_1</ID>219 </input>
<input>
<ID>SEL_2</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>449</ID>
<type>GA_LED</type>
<position>14,122</position>
<input>
<ID>N_in3</ID>221 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>450</ID>
<type>GA_LED</type>
<position>21,122</position>
<input>
<ID>N_in3</ID>222 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>451</ID>
<type>GA_LED</type>
<position>28,122</position>
<input>
<ID>N_in3</ID>223 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>452</ID>
<type>AA_LABEL</type>
<position>13.5,120</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>453</ID>
<type>AA_LABEL</type>
<position>20.5,120</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>454</ID>
<type>AA_LABEL</type>
<position>28,120</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>455</ID>
<type>AA_LABEL</type>
<position>28,118</position>
<gparam>LABEL_TEXT A>B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>AA_LABEL</type>
<position>13.5,118</position>
<gparam>LABEL_TEXT AB</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>457</ID>
<type>AA_LABEL</type>
<position>20.5,118</position>
<gparam>LABEL_TEXT A=B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>AA_AND2</type>
<position>146,55.5</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>459</ID>
<type>AE_OR2</type>
<position>146,60</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>AI_XOR2</type>
<position>146.5,64.5</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>461</ID>
<type>AA_AND2</type>
<position>145.5,32.5</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_OR2</type>
<position>145.5,37</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>463</ID>
<type>AI_XOR2</type>
<position>146,41.5</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>464</ID>
<type>AI_XOR2</type>
<position>78,80</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>465</ID>
<type>AA_AND2</type>
<position>69,68.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>466</ID>
<type>AE_SMALL_INVERTER</type>
<position>61.5,67.5</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>467</ID>
<type>AI_XOR2</type>
<position>71.5,56</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>468</ID>
<type>AA_AND2</type>
<position>68.5,46</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>191 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>469</ID>
<type>AE_SMALL_INVERTER</type>
<position>60,45</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>470</ID>
<type>AI_XOR2</type>
<position>95,60.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>471</ID>
<type>AA_AND2</type>
<position>102.5,52</position>
<input>
<ID>IN_0</ID>196 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>472</ID>
<type>AE_SMALL_INVERTER</type>
<position>95.5,53</position>
<input>
<ID>IN_0</ID>194 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>473</ID>
<type>AE_OR2</type>
<position>121,46</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>478</ID>
<type>AA_LABEL</type>
<position>76,91.5</position>
<gparam>LABEL_TEXT 2 bit Substraction</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>489</ID>
<type>AI_XOR2</type>
<position>63,26</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>490</ID>
<type>AA_AND2</type>
<position>45,2</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>491</ID>
<type>AI_XOR2</type>
<position>73,17</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>492</ID>
<type>AA_AND2</type>
<position>71.5,-6.5</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>493</ID>
<type>AI_XOR2</type>
<position>101.5,16</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_AND2</type>
<position>101.5,3</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>AE_OR2</type>
<position>113,-5.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>496</ID>
<type>AA_LABEL</type>
<position>77.5,34.5</position>
<gparam>LABEL_TEXT 2 bit Addition</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>504</ID>
<type>AA_TOGGLE</type>
<position>10.5,107</position>
<output>
<ID>OUT_0</ID>193 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>505</ID>
<type>AA_TOGGLE</type>
<position>15,107</position>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_TOGGLE</type>
<position>19.5,107</position>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>507</ID>
<type>AA_TOGGLE</type>
<position>23,107</position>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>508</ID>
<type>AA_TOGGLE</type>
<position>28,107</position>
<output>
<ID>OUT_0</ID>220 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_TOGGLE</type>
<position>31,107</position>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>510</ID>
<type>AA_TOGGLE</type>
<position>34,107</position>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_LABEL</type>
<position>11.5,109.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>512</ID>
<type>AA_LABEL</type>
<position>15.5,109.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>513</ID>
<type>AA_LABEL</type>
<position>19.5,109.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>514</ID>
<type>AA_LABEL</type>
<position>23.5,109.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>515</ID>
<type>AA_LABEL</type>
<position>31,109.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>516</ID>
<type>AA_LABEL</type>
<position>34.5,109.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>AA_LABEL</type>
<position>28,109.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>535</ID>
<type>AA_AND2</type>
<position>72.5,-33</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>209 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>536</ID>
<type>AA_AND2</type>
<position>91.5,-58.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>537</ID>
<type>AA_AND2</type>
<position>73,-85.5</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>538</ID>
<type>AE_OR2</type>
<position>128.5,-39</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>539</ID>
<type>AE_OR2</type>
<position>132.5,-79.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>541</ID>
<type>FF_GND</type>
<position>159,12</position>
<output>
<ID>OUT_0</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>542</ID>
<type>FF_GND</type>
<position>160,42.5</position>
<output>
<ID>OUT_0</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>544</ID>
<type>FF_GND</type>
<position>159.5,58.5</position>
<output>
<ID>OUT_0</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-84,10.5,105</points>
<connection>
<GID>504</GID>
<name>OUT_0</name></connection>
<intersection>-84 19</intersection>
<intersection>-54 17</intersection>
<intersection>-32 15</intersection>
<intersection>-7.5 13</intersection>
<intersection>18 22</intersection>
<intersection>42.5 11</intersection>
<intersection>45 4</intersection>
<intersection>58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,58.5,67.5,58.5</points>
<intersection>10.5 0</intersection>
<intersection>67.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>10.5,45,58,45</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>67.5,57,67.5,58.5</points>
<intersection>57 28</intersection>
<intersection>58.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>10.5,42.5,143,42.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection>
<intersection>136 23</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>10.5,-7.5,68.5,-7.5</points>
<connection>
<GID>492</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>10.5,-32,69.5,-32</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>10.5,-54,33,-54</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>10.5,-84,42.5,-84</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>10.5,18,70,18</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>136,33.5,136,42.5</points>
<intersection>33.5 26</intersection>
<intersection>38 24</intersection>
<intersection>42.5 11</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>136,38,142.5,38</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>136 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>136,33.5,142.5,33.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>136 23</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>67.5,57,68.5,57</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>67.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,56,83.5,61.5</points>
<intersection>56 2</intersection>
<intersection>61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,61.5,92,61.5</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection>
<intersection>87 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,56,83.5,56</points>
<connection>
<GID>467</GID>
<name>OUT</name></connection>
<intersection>83.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>87,53,87,61.5</points>
<intersection>53 4</intersection>
<intersection>61.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>87,53,93.5,53</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>87 3</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,45,93,46</points>
<intersection>45 1</intersection>
<intersection>46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,45,118,45</points>
<connection>
<GID>473</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,46,93,46</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97.5,53,99.5,53</points>
<connection>
<GID>472</GID>
<name>OUT_0</name></connection>
<connection>
<GID>471</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,51,43.5,64.5</points>
<intersection>51 1</intersection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,51,99.5,51</points>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection>
<intersection>91 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,64.5,72.5,64.5</points>
<intersection>43.5 0</intersection>
<intersection>72.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72.5,64.5,72.5,68.5</points>
<intersection>64.5 2</intersection>
<intersection>68.5 7</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>91,51,91,59.5</points>
<intersection>51 1</intersection>
<intersection>59.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>91,59.5,92,59.5</points>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>91 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>72,68.5,72.5,68.5</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<intersection>72.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,47,110.5,52</points>
<intersection>47 1</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,47,118,47</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,52,110.5,52</points>
<connection>
<GID>471</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,17,98.5,17</points>
<connection>
<GID>491</GID>
<name>OUT</name></connection>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>82.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>82.5,4,82.5,17</points>
<intersection>4 10</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>82.5,4,98.5,4</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>82.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-6.5,110,-6.5</points>
<connection>
<GID>492</GID>
<name>OUT</name></connection>
<connection>
<GID>495</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,2,98.5,2</points>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<connection>
<GID>490</GID>
<name>OUT</name></connection>
<intersection>97.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>97.5,2,97.5,15</points>
<intersection>2 1</intersection>
<intersection>15 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>97.5,15,98.5,15</points>
<connection>
<GID>493</GID>
<name>IN_1</name></connection>
<intersection>97.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-4.5,106.5,3</points>
<intersection>-4.5 6</intersection>
<intersection>3 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>106.5,-4.5,110,-4.5</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>104.5,3,106.5,3</points>
<connection>
<GID>494</GID>
<name>OUT</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-38,85,-33</points>
<intersection>-38 1</intersection>
<intersection>-33 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-38,125.5,-38</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>75.5,-33,85,-33</points>
<connection>
<GID>535</GID>
<name>OUT</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>95,-78.5,95,-71</points>
<intersection>-78.5 4</intersection>
<intersection>-71 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>95,-78.5,129.5,-78.5</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>92.5,-71,95,-71</points>
<connection>
<GID>444</GID>
<name>OUT</name></connection>
<intersection>95 3</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-85.5,88,-80.5</points>
<intersection>-85.5 4</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-80.5,129.5,-80.5</points>
<connection>
<GID>539</GID>
<name>IN_1</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>76,-85.5,88,-85.5</points>
<connection>
<GID>537</GID>
<name>OUT</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-40,125.5,-40</points>
<connection>
<GID>538</GID>
<name>IN_1</name></connection>
<intersection>109 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>109,-46.5,109,-40</points>
<intersection>-46.5 12</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>93,-46.5,109,-46.5</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<intersection>109 9</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-72,76.5,-47.5</points>
<intersection>-72 16</intersection>
<intersection>-57.5 6</intersection>
<intersection>-54.5 13</intersection>
<intersection>-47.5 15</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>76.5,-57.5,88.5,-57.5</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>48.5,-54.5,76.5,-54.5</points>
<intersection>48.5 17</intersection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>76.5,-47.5,87,-47.5</points>
<connection>
<GID>442</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>76.5,-72,86.5,-72</points>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>48.5,-55.5,48.5,-54.5</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<intersection>-54.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,-79.5,161.5,-79.5</points>
<connection>
<GID>539</GID>
<name>OUT</name></connection>
<intersection>161.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>161.5,-79.5,161.5,11</points>
<connection>
<GID>446</GID>
<name>IN_2</name></connection>
<intersection>-79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-37,47.5,-37</points>
<connection>
<GID>436</GID>
<name>OUT_0</name></connection>
<intersection>47.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>47.5,-37,47.5,-34</points>
<intersection>-37 1</intersection>
<intersection>-34 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>47.5,-34,69.5,-34</points>
<connection>
<GID>535</GID>
<name>IN_1</name></connection>
<intersection>47.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-84.5,51,-84</points>
<intersection>-84.5 1</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-84.5,70,-84.5</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-84,51,-84</points>
<connection>
<GID>434</GID>
<name>OUT_0</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-48,60.5,-42</points>
<intersection>-48 4</intersection>
<intersection>-42 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60.5,-42,68.5,-42</points>
<connection>
<GID>441</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47,-48,60.5,-48</points>
<connection>
<GID>433</GID>
<name>OUT_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-77.5,50.5,-73</points>
<intersection>-77.5 4</intersection>
<intersection>-73 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,-73,50.5,-73</points>
<connection>
<GID>435</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-77.5,68,-77.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-55.5,42.5,-55.5</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>39 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>39,-55.5,39,-55</points>
<connection>
<GID>437</GID>
<name>OUT</name></connection>
<intersection>-55.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>39,-61.5,43,-61.5</points>
<connection>
<GID>439</GID>
<name>OUT</name></connection>
<connection>
<GID>440</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-61.5,75,-59.5</points>
<intersection>-61.5 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-59.5,88.5,-59.5</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-61.5,75,-61.5</points>
<connection>
<GID>440</GID>
<name>OUT_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-41,87,-41</points>
<connection>
<GID>441</GID>
<name>OUT</name></connection>
<intersection>87 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>87,-45.5,87,-41</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-70,86.5,-70</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>74 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>74,-78.5,74,-70</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<intersection>-70 1</intersection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,15,165.5,101</points>
<connection>
<GID>446</GID>
<name>SEL_0</name></connection>
<connection>
<GID>447</GID>
<name>SEL_0</name></connection>
<connection>
<GID>448</GID>
<name>SEL_0</name></connection>
<intersection>101 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>34,101,34,105</points>
<connection>
<GID>510</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34,101,165.5,101</points>
<intersection>34 1</intersection>
<intersection>165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,15,164.5,98.5</points>
<connection>
<GID>446</GID>
<name>SEL_1</name></connection>
<connection>
<GID>447</GID>
<name>SEL_1</name></connection>
<connection>
<GID>448</GID>
<name>SEL_1</name></connection>
<intersection>98.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,98.5,31,105</points>
<connection>
<GID>509</GID>
<name>OUT_0</name></connection>
<intersection>98.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31,98.5,164.5,98.5</points>
<intersection>31 1</intersection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,45.5,163.5,96.5</points>
<connection>
<GID>447</GID>
<name>SEL_2</name></connection>
<connection>
<GID>448</GID>
<name>SEL_2</name></connection>
<intersection>96.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>28,96.5,28,105</points>
<connection>
<GID>508</GID>
<name>OUT_0</name></connection>
<intersection>96.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28,96.5,163.5,96.5</points>
<intersection>28 1</intersection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,123,14,140.5</points>
<connection>
<GID>449</GID>
<name>N_in3</name></connection>
<intersection>140.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,140.5,185,140.5</points>
<intersection>14 0</intersection>
<intersection>185 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>185,10,185,140.5</points>
<intersection>10 3</intersection>
<intersection>140.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>167.5,10,185,10</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<intersection>185 2</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,130,182.5,130</points>
<intersection>21 3</intersection>
<intersection>182.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21,123,21,130</points>
<connection>
<GID>450</GID>
<name>N_in3</name></connection>
<intersection>130 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>182.5,40,182.5,130</points>
<intersection>40 5</intersection>
<intersection>130 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>167.5,40,182.5,40</points>
<connection>
<GID>447</GID>
<name>OUT</name></connection>
<intersection>182.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,126.5,176.5,126.5</points>
<intersection>28 7</intersection>
<intersection>176.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>176.5,56,176.5,126.5</points>
<intersection>56 4</intersection>
<intersection>126.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>167.5,56,176.5,56</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>176.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>28,123,28,126.5</points>
<connection>
<GID>451</GID>
<name>N_in3</name></connection>
<intersection>126.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,36.5,152,60.5</points>
<intersection>36.5 2</intersection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,60.5,152,60.5</points>
<connection>
<GID>470</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,36.5,161.5,36.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,7,145,46</points>
<intersection>7 2</intersection>
<intersection>46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,46,145,46</points>
<connection>
<GID>473</GID>
<name>OUT</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145,7,161.5,7</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,26,153.5,53.5</points>
<intersection>26 1</intersection>
<intersection>53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,26,153.5,26</points>
<connection>
<GID>489</GID>
<name>OUT</name></connection>
<intersection>153.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153.5,53.5,161.5,53.5</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>153.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,16,154.5,37.5</points>
<intersection>16 2</intersection>
<intersection>37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154.5,37.5,161.5,37.5</points>
<connection>
<GID>447</GID>
<name>IN_1</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,16,154.5,16</points>
<connection>
<GID>493</GID>
<name>OUT</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-5.5,154.5,9</points>
<intersection>-5.5 2</intersection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154.5,9,161.5,9</points>
<connection>
<GID>446</GID>
<name>IN_1</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-5.5,154.5,-5.5</points>
<connection>
<GID>495</GID>
<name>OUT</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-39,153,54.5</points>
<intersection>-39 1</intersection>
<intersection>54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-39,153,-39</points>
<connection>
<GID>538</GID>
<name>OUT</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153,54.5,161.5,54.5</points>
<connection>
<GID>448</GID>
<name>IN_2</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-58.5,151,38</points>
<intersection>-58.5 2</intersection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,38,161.5,38</points>
<intersection>151 0</intersection>
<intersection>161.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-58.5,151,-58.5</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>161.5,38,161.5,38.5</points>
<connection>
<GID>447</GID>
<name>IN_2</name></connection>
<intersection>38 1</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,55.5,161.5,55.5</points>
<connection>
<GID>458</GID>
<name>OUT</name></connection>
<connection>
<GID>448</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,32.5,156,39.5</points>
<intersection>32.5 2</intersection>
<intersection>39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,39.5,161.5,39.5</points>
<connection>
<GID>447</GID>
<name>IN_3</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,32.5,156,32.5</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159,13,161.5,13</points>
<connection>
<GID>541</GID>
<name>OUT_0</name></connection>
<connection>
<GID>446</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160,43.5,161.5,43.5</points>
<connection>
<GID>542</GID>
<name>OUT_0</name></connection>
<connection>
<GID>447</GID>
<name>IN_7</name></connection>
<intersection>161.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>161.5,42.5,161.5,43.5</points>
<connection>
<GID>447</GID>
<name>IN_6</name></connection>
<intersection>43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,58.5,161.5,59.5</points>
<connection>
<GID>448</GID>
<name>IN_6</name></connection>
<connection>
<GID>448</GID>
<name>IN_7</name></connection>
<intersection>59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159.5,59.5,161.5,59.5</points>
<connection>
<GID>544</GID>
<name>OUT_0</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,57.5,155,60</points>
<intersection>57.5 1</intersection>
<intersection>60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155,57.5,161.5,57.5</points>
<connection>
<GID>448</GID>
<name>IN_5</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149,60,155,60</points>
<connection>
<GID>459</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,56.5,155.5,64.5</points>
<intersection>56.5 1</intersection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,56.5,161.5,56.5</points>
<connection>
<GID>448</GID>
<name>IN_4</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149.5,64.5,155.5,64.5</points>
<connection>
<GID>460</GID>
<name>OUT</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,37,150,40</points>
<intersection>37 2</intersection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,40,158.5,40</points>
<intersection>150 0</intersection>
<intersection>158.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,37,150,37</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>150 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>158.5,40,158.5,41.5</points>
<intersection>40 1</intersection>
<intersection>41.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>158.5,41.5,161.5,41.5</points>
<connection>
<GID>447</GID>
<name>IN_5</name></connection>
<intersection>158.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,40.5,155,41.5</points>
<intersection>40.5 1</intersection>
<intersection>41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155,40.5,161.5,40.5</points>
<connection>
<GID>447</GID>
<name>IN_4</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149,41.5,155,41.5</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,85,138,85</points>
<intersection>15 3</intersection>
<intersection>73 32</intersection>
<intersection>138 25</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-73,15,105</points>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection>
<intersection>-73 22</intersection>
<intersection>-60.5 20</intersection>
<intersection>-40 18</intersection>
<intersection>1 16</intersection>
<intersection>27 14</intersection>
<intersection>67.5 4</intersection>
<intersection>85 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15,67.5,59.5,67.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>15,27,60,27</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>15,1,42,1</points>
<connection>
<GID>490</GID>
<name>IN_1</name></connection>
<intersection>15 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>15,-40,68.5,-40</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>15,-60.5,33,-60.5</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>15,-73,41,-73</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>138,56.5,138,85</points>
<intersection>56.5 30</intersection>
<intersection>61 28</intersection>
<intersection>65.5 26</intersection>
<intersection>85 1</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>138,65.5,143.5,65.5</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>138 25</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>138,61,143,61</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>138 25</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>138,56.5,143,56.5</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>138 25</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>73,81,73,85</points>
<intersection>81 33</intersection>
<intersection>85 1</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>73,81,75,81</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>73 32</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,74.5,139,74.5</points>
<intersection>23 3</intersection>
<intersection>73 34</intersection>
<intersection>139 24</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-79.5,23,105</points>
<connection>
<GID>507</GID>
<name>OUT_0</name></connection>
<intersection>-79.5 23</intersection>
<intersection>-62.5 21</intersection>
<intersection>-48 19</intersection>
<intersection>3 17</intersection>
<intersection>25 15</intersection>
<intersection>69.5 4</intersection>
<intersection>74.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23,69.5,66,69.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>23,25,60,25</points>
<connection>
<GID>489</GID>
<name>IN_1</name></connection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>23,3,42,3</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>23,-48,41,-48</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>23,-62.5,33,-62.5</points>
<connection>
<GID>439</GID>
<name>IN_1</name></connection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>23,-79.5,68,-79.5</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>139,54.5,139,74.5</points>
<intersection>54.5 32</intersection>
<intersection>59 30</intersection>
<intersection>63.5 27</intersection>
<intersection>74.5 1</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>139,63.5,143.5,63.5</points>
<connection>
<GID>460</GID>
<name>IN_1</name></connection>
<intersection>139 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>139,59,143,59</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<intersection>139 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>139,54.5,143,54.5</points>
<connection>
<GID>458</GID>
<name>IN_1</name></connection>
<intersection>139 24</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>73,74.5,73,79</points>
<intersection>74.5 1</intersection>
<intersection>79 35</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>73,79,75,79</points>
<connection>
<GID>464</GID>
<name>IN_1</name></connection>
<intersection>73 34</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>63.5,67.5,66,67.5</points>
<connection>
<GID>466</GID>
<name>OUT_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,55,68.5,55</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<intersection>19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19.5,-86.5,19.5,105</points>
<connection>
<GID>506</GID>
<name>OUT_0</name></connection>
<intersection>-86.5 18</intersection>
<intersection>-56 16</intersection>
<intersection>-37 14</intersection>
<intersection>-5.5 12</intersection>
<intersection>16 10</intersection>
<intersection>40.5 20</intersection>
<intersection>47 4</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19.5,47,65.5,47</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>19.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>19.5,16,70,16</points>
<connection>
<GID>491</GID>
<name>IN_1</name></connection>
<intersection>19.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>19.5,-5.5,68.5,-5.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>19.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>19.5,-37,38,-37</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<intersection>19.5 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>19.5,-56,33,-56</points>
<connection>
<GID>437</GID>
<name>IN_1</name></connection>
<intersection>19.5 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>19.5,-86.5,70,-86.5</points>
<connection>
<GID>537</GID>
<name>IN_1</name></connection>
<intersection>19.5 3</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>19.5,40.5,143,40.5</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<intersection>19.5 3</intersection>
<intersection>137 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>137,31.5,137,40.5</points>
<intersection>31.5 25</intersection>
<intersection>36 22</intersection>
<intersection>40.5 20</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>137,36,142.5,36</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<intersection>137 21</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>137,31.5,142.5,31.5</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<intersection>137 21</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,45,65.5,45</points>
<connection>
<GID>469</GID>
<name>OUT_0</name></connection>
<connection>
<GID>468</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,52.5,120,80</points>
<intersection>52.5 13</intersection>
<intersection>80 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>81,80,120,80</points>
<connection>
<GID>464</GID>
<name>OUT</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>120,52.5,161.5,52.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-6.00815e-006,0,44.2,-46.2</PageViewport></page 5>
<page 6>
<PageViewport>-6.00815e-006,0,44.2,-46.2</PageViewport></page 6>
<page 7>
<PageViewport>-6.00815e-006,0,44.2,-46.2</PageViewport></page 7>
<page 8>
<PageViewport>-6.00815e-006,0,44.2,-46.2</PageViewport></page 8>
<page 9>
<PageViewport>-6.00815e-006,0,44.2,-46.2</PageViewport></page 9></circuit>